module pscontroller(CLOCK_50, resetn, ps2_clk, ps2_keyboard_data);

	//Input
	input CLOCK_50;
	input resetn;
		
	
	//Output
	
	//Wire

endmodule