`default_nettype none
`include "params.vh"

module vga_adapter(
    resetn, clock, color, x, y, write,
    VGA_R, VGA_G, VGA_B, VGA_HS, VGA_VS, VGA_BLANK_N, VGA_SYNC_N, VGA_CLK,
    player_tile_x, player_tile_y, player_dir
);

    // The VGA resolution, which can be set to "640x480", "320x240", and "160x120"
    parameter RESOLUTION = "640x480";

    // 3 bits per R/G/B = 9-bit color
    parameter COLOR_DEPTH = 9;

    // Number of VGA pixel X coordinate (column) and Y coordinate (row) bits
    parameter nX = (RESOLUTION == "640x480") ? 10 :
                   ((RESOLUTION == "320x240") ? 9 : 8);
    parameter nY = (RESOLUTION == "640x480") ? 9  :
                   ((RESOLUTION == "320x240") ? 8 : 7);

    // Number of address bits on the video memory
    parameter Mn = (RESOLUTION == "640x480") ? 19 :
                   ((RESOLUTION == "320x240") ? 17 : 15);

    // Number of columns and rows in the video memory
    parameter COLS = (RESOLUTION == "640x480") ? 640 :
                     ((RESOLUTION == "320x240") ? 320 : 160);
    parameter ROWS = (RESOLUTION == "640x480") ? 480 :
                     ((RESOLUTION == "320x240") ? 240 : 120);

    input  wire                        resetn;
    input  wire                        clock;
	 
	     // Player tile position (grid 0..29 × 0..11) and direction
    input  wire [4:0] player_tile_x;
    input  wire [4:0] player_tile_y;
    input  wire [1:0] player_dir;


    // These are *not* used now – background comes from ROM
    input  wire [COLOR_DEPTH-1:0]      color;
    input  wire [nX-1:0]               x;
    input  wire [nY-1:0]               y;
    input  wire                        write;

    output wire [7:0]                  VGA_R;
    output wire [7:0]                  VGA_G;
    output wire [7:0]                  VGA_B;
    output wire                        VGA_HS;
    output wire                        VGA_VS;
    output wire                        VGA_BLANK_N;
    output wire                        VGA_SYNC_N;
    output wire                        VGA_CLK;

    // ----------------------------------------------------------------
    // Local signals
    // ----------------------------------------------------------------
    reg         clock_25;   // 25 MHz derived from 50 MHz
    wire [Mn-1:0] controller_to_video_memory_addr;
    wire [COLOR_DEPTH-1:0] rom_color;

	 

	

    // ----------------------------------------------------------------
    // 50 MHz -> 25 MHz clock divider (replaces vga_pll)
    // ----------------------------------------------------------------
    always @(posedge clock or negedge resetn) begin
        if (!resetn)
            clock_25 <= 1'b0;
        else
            clock_25 <= ~clock_25;
    end

    // ----------------------------------------------------------------
    // Background ROM (generated by MegaWizard)
    //   - Make sure *background_rom.v* (not only background_rom_bb.v)
    //     is added to your Quartus project.
    //   - Data width must be 9 bits to match COLOR_DEPTH.
    // ----------------------------------------------------------------
    background_rom VideoMemory (
        .address (controller_to_video_memory_addr),  // which pixel
        .clock   (clock_25),                         // 25 MHz
        .q       (rom_color)                         // 9-bit color
    );

    // ----------------------------------------------------------------
    // VGA Controller: reads ROM, overlays maze from play_map.v
    // ----------------------------------------------------------------
	 
    /*vga_controller controller(
        .vga_clock      (clock_25),
        .resetn         (resetn),
        .pixel_color    (rom_color),
        .memory_address (controller_to_video_memory_addr),
        .VGA_R          (VGA_R),
        .VGA_G          (VGA_G),
        .VGA_B          (VGA_B),
        .VGA_HS         (VGA_HS),
        .VGA_VS         (VGA_VS),
        .VGA_BLANK_N    (VGA_BLANK_N),
        .VGA_SYNC_N     (VGA_SYNC_N),
        .VGA_CLK        (VGA_CLK),
        .player_x       (player_x),
        .player_y       (player_y)
    );
	 */
	 
    vga_controller controller(
        .vga_clock      (clock_25),
        .resetn         (resetn),
        .pixel_color    (rom_color),
        .memory_address (controller_to_video_memory_addr),
        .VGA_R          (VGA_R),
        .VGA_G          (VGA_G),
        .VGA_B          (VGA_B),
        .VGA_HS         (VGA_HS),
        .VGA_VS         (VGA_VS),
        .VGA_BLANK_N    (VGA_BLANK_N),
        .VGA_SYNC_N     (VGA_SYNC_N),
        .VGA_CLK        (VGA_CLK),
        .player_x       (player_tile_x),
        .player_y       (player_tile_y),
        .player_dir     (player_dir)
    );

	 
    defparam controller.RESOLUTION  = RESOLUTION;
    defparam controller.COLOR_DEPTH = COLOR_DEPTH;
    defparam controller.nX          = nX;
    defparam controller.nY          = nY;
    defparam controller.Mn          = Mn;
    defparam controller.ROWS        = ROWS;
    defparam controller.COLS        = COLS;

endmodule
