`ifndef PARAMS_VH
`define PARAMS_VH

    `define MAP_WIDTH   21
    `define MAP_HEIGHT  11
    `define DATA_WIDTH  8
    `define ADDR_WIDTH  10

`endif // PARAMS_VH