`ifndef PARAMS_VH
`define PARAMS_VH

    `define MAP_WIDTH   30        // 30 columns
    `define MAP_HEIGHT  12        // 12 rows

    `define DATA_WIDTH  8
    `define ADDR_WIDTH  10

`endif // PARAMS_VH
